entity ieee;

